module Clock (
    input [0:0] clk,
    output [0:0] uart_clk_16
);


    
endmodule