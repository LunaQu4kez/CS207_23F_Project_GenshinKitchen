module Automatic (
    input [0:0] clk,
    input [7:0] out_bits,
    input [0:0] out_valid,
    input [0:0] in_ready,
    input [0:0] mode,
    input [15:0] script,
    output [7:0] pc,
    output [7:0] in_bits
);

    

    
endmodule