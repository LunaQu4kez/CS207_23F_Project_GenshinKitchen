`timescale 1ns / 1ps

module Top(
    input [4:0] button,
    input [7:0] switches,

    output [7:0] led,
    output [7:0] led2,
    
    input clk,
    input rx,
    output tx
);

    wire uart_clk_16;
        
    reg [7:0] dataIn_bits;
    wire dataIn_ready;
    reg state_flag = 1'b0; // 0 not start, 1 start
    
    wire [7:0] dataOut_bits;
    wire dataOut_valid;
    
    wire script_mode;
    wire [7:0] pc;
    wire [15:0] script;


    ScriptMem script_mem_module(
        .clock(uart_clk_16),   // please use the same clock as UART module
        .reset(0),           // please use the same reset as UART module
    
        .dataOut_bits(dataOut_bits), // please connect to io_dataOut_bits of UART module
        .dataOut_valid(dataOut_valid), // please connect to io_dataOut_valid of UART module
    
        .script_mode(script_mode), // output 1 when loading script from UART.
                                   // at this time, you should not use dataOut_bits or use pc and script.
    
        .pc(pc), // (a) give a program counter (address) to ScriptMem.
        .script(script) // referring (a), returning the corresponding instructions of pc
    );

    UART uart_module(
        .clock(uart_clk_16),     // uart clock. Please use 16 x BultRate. (e.g. 9600 * 16 = 153600Hz)
        .reset(0),               // reset
  
        .io_pair_rx(rx),          // rx, connect to R5 please
        .io_pair_tx(tx),         // tx, connect to T4 please
        
        .io_dataIn_bits(dataIn_bits),     // (a) byte from DevelopmentBoard => GenshinKitchen
        .io_dataIn_ready(dataIn_ready),   // referring (a) pulse 1 after a byte tramsmit success.
        
        .io_dataOut_bits(dataOut_bits),     // (b) byte from GenshinKitchen => DevelopmentBoard, only available if io_dataOut_valid=1
        .io_dataOut_valid(dataOut_valid)  // referring (b)
    );

    Clock clock(
        .clk(clk),
        .uart_clk_16(uart_clk_16)
    );

    always @(posedge uart_clk_16) begin
        if (dataIn_ready) begin
            if (switches[7] & ~state_flag) begin
                state_flag <= 1'b1;
                dataIn_bits <= 8'b0000_0101;
            end
            else if (~switches[7] & state_flag) begin
                state_flag <= 1'b0;
                dataIn_bits <= 8'b0000_1001;
            end
        end
        else begin
            dataIn_bits <= 8'b0000_0000;
        end
    end




endmodule